module ScoreDisplay();
endmodule